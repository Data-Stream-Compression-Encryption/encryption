module S_Box_1(in, out);
  input [5:0] in;
  output [3:0] out;
  
endmodule
