`timescale 1 ns/ 1 ps

module S_Box_1(in, out);
  input [5:0] in;
  output [3:0] out;
  
  assign out =  (in == 6'b000000) ? 4'd14 :
                (in == 6'b000010) ? 4'd4  :
                (in == 6'b000100) ? 4'd13 :
                (in == 6'b000110) ? 4'd1  :
                (in == 6'b001000) ? 4'd2  :
                (in == 6'b001010) ? 4'd15 :
                (in == 6'b001100) ? 4'd11 :
                (in == 6'b001110) ? 4'd8  :
                (in == 6'b010000) ? 4'd3  :
                (in == 6'b010010) ? 4'd10 :
                (in == 6'b010100) ? 4'd6  :
                (in == 6'b010110) ? 4'd12 :
                (in == 6'b011000) ? 4'd5  :
                (in == 6'b011010) ? 4'd9  :
                (in == 6'b011100) ? 4'd0  :
                (in == 6'b011110) ? 4'd7  :
                
                (in == 6'b000001) ? 4'd0  :
                (in == 6'b000011) ? 4'd15 :
                (in == 6'b000101) ? 4'd7  :
                (in == 6'b000111) ? 4'd4  :
                (in == 6'b001001) ? 4'd14 :
                (in == 6'b001011) ? 4'd2  :
                (in == 6'b001101) ? 4'd13 :
                (in == 6'b001111) ? 4'd1  :
                (in == 6'b010001) ? 4'd10 :
                (in == 6'b010011) ? 4'd6  :
                (in == 6'b010101) ? 4'd12 :
                (in == 6'b010111) ? 4'd11 :
                (in == 6'b011001) ? 4'd9  :
                (in == 6'b011011) ? 4'd5  :
                (in == 6'b011101) ? 4'd3  :
                (in == 6'b011111) ? 4'd8  :
                
                (in == 6'b100000) ? 4'd4  :
                (in == 6'b100010) ? 4'd1  :
                (in == 6'b100100) ? 4'd14 :
                (in == 6'b100110) ? 4'd8  :
                (in == 6'b101000) ? 4'd13 :
                (in == 6'b101010) ? 4'd6  :
                (in == 6'b101100) ? 4'd2  :
                (in == 6'b101110) ? 4'd11 :
                (in == 6'b110000) ? 4'd15 :
                (in == 6'b110010) ? 4'd12 :
                (in == 6'b110100) ? 4'd9  :
                (in == 6'b110110) ? 4'd7  :
                (in == 6'b111000) ? 4'd3  :
                (in == 6'b111010) ? 4'd10 :
                (in == 6'b111100) ? 4'd5  :
                (in == 6'b111110) ? 4'd0  :
                
                (in == 6'b100001) ? 4'd15 :
                (in == 6'b100011) ? 4'd12 :
                (in == 6'b100101) ? 4'd8  :
                (in == 6'b100111) ? 4'd2  :
                (in == 6'b101001) ? 4'd4  :
                (in == 6'b101011) ? 4'd9  :
                (in == 6'b101101) ? 4'd1  :
                (in == 6'b101111) ? 4'd7  :
                (in == 6'b110001) ? 4'd5  :
                (in == 6'b110011) ? 4'd11 :
                (in == 6'b110101) ? 4'd3  :
                (in == 6'b110111) ? 4'd14 :
                (in == 6'b111001) ? 4'd10 :
                (in == 6'b111011) ? 4'd0  :
                (in == 6'b111101) ? 4'd6  : 4'd13; 
  
endmodule
