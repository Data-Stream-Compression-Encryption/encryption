/*

Module:   TB_DES
Purpose:  Tests the DES Algorithm in accordance with the procedure described at
          http://people.csail.mit.edu/rivest/pubs/Riv85.txt

*/

`timescale 1 ns/ 1 ps

module TB_DES;
  
  reg clk;
  reg [63:0] in;
  reg [63:0] out;
  
  
endmodule